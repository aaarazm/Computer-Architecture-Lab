module EX(
	PC_In,
	Signed_EX_imm_24,
	Branch_Address
);

input[31:0] PC_In;
input[23:0] Signed_EX_imm_24;
output [31:0]Branch_Address;

endmodule 
