module helloWorld(
    a, b, w
);
    input a, b;
    output w;
    assign w = a || b;
endmodule