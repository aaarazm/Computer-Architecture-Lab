module ARM(clk);
    input clk;
    IF IF_inst(

    );

endmodule